library verilog;
use verilog.vl_types.all;
entity DigChoose_vlg_vec_tst is
end DigChoose_vlg_vec_tst;
