library verilog;
use verilog.vl_types.all;
entity ioRead_test is
end ioRead_test;
