library verilog;
use verilog.vl_types.all;
entity showall_test is
end showall_test;
